VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1050.310 BY 1061.030 ;
  PIN iClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END iClk
  PIN iRst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END iRst_n
  PIN iSDAT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END iSDAT
  PIN iSVAL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END iSVAL
  PIN iSize[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END iSize[0]
  PIN iSize[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 1057.030 875.290 1061.030 ;
    END
  END iSize[1]
  PIN iSize[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 0.000 975.110 4.000 ;
    END
  END iSize[2]
  PIN iValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END iValid
  PIN oSDAT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 1057.030 525.230 1061.030 ;
    END
  END oSDAT
  PIN oSVAL
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 1057.030 175.170 1061.030 ;
    END
  END oSVAL
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1050.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1050.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1050.160 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 1045.785 1044.850 1048.615 ;
        RECT 5.330 1040.345 1044.850 1043.175 ;
        RECT 5.330 1034.905 1044.850 1037.735 ;
        RECT 5.330 1029.465 1044.850 1032.295 ;
        RECT 5.330 1024.025 1044.850 1026.855 ;
        RECT 5.330 1018.585 1044.850 1021.415 ;
        RECT 5.330 1013.145 1044.850 1015.975 ;
        RECT 5.330 1007.705 1044.850 1010.535 ;
        RECT 5.330 1002.265 1044.850 1005.095 ;
        RECT 5.330 996.825 1044.850 999.655 ;
        RECT 5.330 991.385 1044.850 994.215 ;
        RECT 5.330 985.945 1044.850 988.775 ;
        RECT 5.330 980.505 1044.850 983.335 ;
        RECT 5.330 975.065 1044.850 977.895 ;
        RECT 5.330 969.625 1044.850 972.455 ;
        RECT 5.330 964.185 1044.850 967.015 ;
        RECT 5.330 958.745 1044.850 961.575 ;
        RECT 5.330 953.305 1044.850 956.135 ;
        RECT 5.330 947.865 1044.850 950.695 ;
        RECT 5.330 942.425 1044.850 945.255 ;
        RECT 5.330 936.985 1044.850 939.815 ;
        RECT 5.330 931.545 1044.850 934.375 ;
        RECT 5.330 926.105 1044.850 928.935 ;
        RECT 5.330 920.665 1044.850 923.495 ;
        RECT 5.330 915.225 1044.850 918.055 ;
        RECT 5.330 909.785 1044.850 912.615 ;
        RECT 5.330 904.345 1044.850 907.175 ;
        RECT 5.330 898.905 1044.850 901.735 ;
        RECT 5.330 893.465 1044.850 896.295 ;
        RECT 5.330 888.025 1044.850 890.855 ;
        RECT 5.330 882.585 1044.850 885.415 ;
        RECT 5.330 877.145 1044.850 879.975 ;
        RECT 5.330 871.705 1044.850 874.535 ;
        RECT 5.330 866.265 1044.850 869.095 ;
        RECT 5.330 860.825 1044.850 863.655 ;
        RECT 5.330 855.385 1044.850 858.215 ;
        RECT 5.330 849.945 1044.850 852.775 ;
        RECT 5.330 844.505 1044.850 847.335 ;
        RECT 5.330 839.065 1044.850 841.895 ;
        RECT 5.330 833.625 1044.850 836.455 ;
        RECT 5.330 828.185 1044.850 831.015 ;
        RECT 5.330 822.745 1044.850 825.575 ;
        RECT 5.330 817.305 1044.850 820.135 ;
        RECT 5.330 811.865 1044.850 814.695 ;
        RECT 5.330 806.425 1044.850 809.255 ;
        RECT 5.330 800.985 1044.850 803.815 ;
        RECT 5.330 795.545 1044.850 798.375 ;
        RECT 5.330 790.105 1044.850 792.935 ;
        RECT 5.330 784.665 1044.850 787.495 ;
        RECT 5.330 779.225 1044.850 782.055 ;
        RECT 5.330 773.785 1044.850 776.615 ;
        RECT 5.330 768.345 1044.850 771.175 ;
        RECT 5.330 762.905 1044.850 765.735 ;
        RECT 5.330 757.465 1044.850 760.295 ;
        RECT 5.330 752.025 1044.850 754.855 ;
        RECT 5.330 746.585 1044.850 749.415 ;
        RECT 5.330 741.145 1044.850 743.975 ;
        RECT 5.330 735.705 1044.850 738.535 ;
        RECT 5.330 730.265 1044.850 733.095 ;
        RECT 5.330 724.825 1044.850 727.655 ;
        RECT 5.330 719.385 1044.850 722.215 ;
        RECT 5.330 713.945 1044.850 716.775 ;
        RECT 5.330 708.505 1044.850 711.335 ;
        RECT 5.330 703.065 1044.850 705.895 ;
        RECT 5.330 697.625 1044.850 700.455 ;
        RECT 5.330 692.185 1044.850 695.015 ;
        RECT 5.330 686.745 1044.850 689.575 ;
        RECT 5.330 681.305 1044.850 684.135 ;
        RECT 5.330 675.865 1044.850 678.695 ;
        RECT 5.330 670.425 1044.850 673.255 ;
        RECT 5.330 664.985 1044.850 667.815 ;
        RECT 5.330 659.545 1044.850 662.375 ;
        RECT 5.330 654.105 1044.850 656.935 ;
        RECT 5.330 648.665 1044.850 651.495 ;
        RECT 5.330 643.225 1044.850 646.055 ;
        RECT 5.330 637.785 1044.850 640.615 ;
        RECT 5.330 632.345 1044.850 635.175 ;
        RECT 5.330 626.905 1044.850 629.735 ;
        RECT 5.330 621.465 1044.850 624.295 ;
        RECT 5.330 616.025 1044.850 618.855 ;
        RECT 5.330 610.585 1044.850 613.415 ;
        RECT 5.330 605.145 1044.850 607.975 ;
        RECT 5.330 599.705 1044.850 602.535 ;
        RECT 5.330 594.265 1044.850 597.095 ;
        RECT 5.330 588.825 1044.850 591.655 ;
        RECT 5.330 583.385 1044.850 586.215 ;
        RECT 5.330 577.945 1044.850 580.775 ;
        RECT 5.330 572.505 1044.850 575.335 ;
        RECT 5.330 567.065 1044.850 569.895 ;
        RECT 5.330 561.625 1044.850 564.455 ;
        RECT 5.330 556.185 1044.850 559.015 ;
        RECT 5.330 550.745 1044.850 553.575 ;
        RECT 5.330 545.305 1044.850 548.135 ;
        RECT 5.330 539.865 1044.850 542.695 ;
        RECT 5.330 534.425 1044.850 537.255 ;
        RECT 5.330 528.985 1044.850 531.815 ;
        RECT 5.330 523.545 1044.850 526.375 ;
        RECT 5.330 518.105 1044.850 520.935 ;
        RECT 5.330 512.665 1044.850 515.495 ;
        RECT 5.330 507.225 1044.850 510.055 ;
        RECT 5.330 501.785 1044.850 504.615 ;
        RECT 5.330 496.345 1044.850 499.175 ;
        RECT 5.330 490.905 1044.850 493.735 ;
        RECT 5.330 485.465 1044.850 488.295 ;
        RECT 5.330 480.025 1044.850 482.855 ;
        RECT 5.330 474.585 1044.850 477.415 ;
        RECT 5.330 469.145 1044.850 471.975 ;
        RECT 5.330 463.705 1044.850 466.535 ;
        RECT 5.330 458.265 1044.850 461.095 ;
        RECT 5.330 452.825 1044.850 455.655 ;
        RECT 5.330 447.385 1044.850 450.215 ;
        RECT 5.330 441.945 1044.850 444.775 ;
        RECT 5.330 436.505 1044.850 439.335 ;
        RECT 5.330 431.065 1044.850 433.895 ;
        RECT 5.330 425.625 1044.850 428.455 ;
        RECT 5.330 420.185 1044.850 423.015 ;
        RECT 5.330 414.745 1044.850 417.575 ;
        RECT 5.330 409.305 1044.850 412.135 ;
        RECT 5.330 403.865 1044.850 406.695 ;
        RECT 5.330 398.425 1044.850 401.255 ;
        RECT 5.330 392.985 1044.850 395.815 ;
        RECT 5.330 387.545 1044.850 390.375 ;
        RECT 5.330 382.105 1044.850 384.935 ;
        RECT 5.330 376.665 1044.850 379.495 ;
        RECT 5.330 371.225 1044.850 374.055 ;
        RECT 5.330 365.785 1044.850 368.615 ;
        RECT 5.330 360.345 1044.850 363.175 ;
        RECT 5.330 354.905 1044.850 357.735 ;
        RECT 5.330 349.465 1044.850 352.295 ;
        RECT 5.330 344.025 1044.850 346.855 ;
        RECT 5.330 338.585 1044.850 341.415 ;
        RECT 5.330 333.145 1044.850 335.975 ;
        RECT 5.330 327.705 1044.850 330.535 ;
        RECT 5.330 322.265 1044.850 325.095 ;
        RECT 5.330 316.825 1044.850 319.655 ;
        RECT 5.330 311.385 1044.850 314.215 ;
        RECT 5.330 305.945 1044.850 308.775 ;
        RECT 5.330 300.505 1044.850 303.335 ;
        RECT 5.330 295.065 1044.850 297.895 ;
        RECT 5.330 289.625 1044.850 292.455 ;
        RECT 5.330 284.185 1044.850 287.015 ;
        RECT 5.330 278.745 1044.850 281.575 ;
        RECT 5.330 273.305 1044.850 276.135 ;
        RECT 5.330 267.865 1044.850 270.695 ;
        RECT 5.330 262.425 1044.850 265.255 ;
        RECT 5.330 256.985 1044.850 259.815 ;
        RECT 5.330 251.545 1044.850 254.375 ;
        RECT 5.330 246.105 1044.850 248.935 ;
        RECT 5.330 240.665 1044.850 243.495 ;
        RECT 5.330 235.225 1044.850 238.055 ;
        RECT 5.330 229.785 1044.850 232.615 ;
        RECT 5.330 224.345 1044.850 227.175 ;
        RECT 5.330 218.905 1044.850 221.735 ;
        RECT 5.330 213.465 1044.850 216.295 ;
        RECT 5.330 208.025 1044.850 210.855 ;
        RECT 5.330 202.585 1044.850 205.415 ;
        RECT 5.330 197.145 1044.850 199.975 ;
        RECT 5.330 191.705 1044.850 194.535 ;
        RECT 5.330 186.265 1044.850 189.095 ;
        RECT 5.330 180.825 1044.850 183.655 ;
        RECT 5.330 175.385 1044.850 178.215 ;
        RECT 5.330 169.945 1044.850 172.775 ;
        RECT 5.330 164.505 1044.850 167.335 ;
        RECT 5.330 159.065 1044.850 161.895 ;
        RECT 5.330 153.625 1044.850 156.455 ;
        RECT 5.330 148.185 1044.850 151.015 ;
        RECT 5.330 142.745 1044.850 145.575 ;
        RECT 5.330 137.305 1044.850 140.135 ;
        RECT 5.330 131.865 1044.850 134.695 ;
        RECT 5.330 126.425 1044.850 129.255 ;
        RECT 5.330 120.985 1044.850 123.815 ;
        RECT 5.330 115.545 1044.850 118.375 ;
        RECT 5.330 110.105 1044.850 112.935 ;
        RECT 5.330 104.665 1044.850 107.495 ;
        RECT 5.330 99.225 1044.850 102.055 ;
        RECT 5.330 93.785 1044.850 96.615 ;
        RECT 5.330 88.345 1044.850 91.175 ;
        RECT 5.330 82.905 1044.850 85.735 ;
        RECT 5.330 77.465 1044.850 80.295 ;
        RECT 5.330 72.025 1044.850 74.855 ;
        RECT 5.330 66.585 1044.850 69.415 ;
        RECT 5.330 61.145 1044.850 63.975 ;
        RECT 5.330 55.705 1044.850 58.535 ;
        RECT 5.330 50.265 1044.850 53.095 ;
        RECT 5.330 44.825 1044.850 47.655 ;
        RECT 5.330 39.385 1044.850 42.215 ;
        RECT 5.330 33.945 1044.850 36.775 ;
        RECT 5.330 28.505 1044.850 31.335 ;
        RECT 5.330 23.065 1044.850 25.895 ;
        RECT 5.330 17.625 1044.850 20.455 ;
        RECT 5.330 12.185 1044.850 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1044.660 1050.005 ;
      LAYER met1 ;
        RECT 5.520 10.640 1044.660 1050.160 ;
      LAYER met2 ;
        RECT 15.740 1056.750 174.610 1057.810 ;
        RECT 175.450 1056.750 524.670 1057.810 ;
        RECT 525.510 1056.750 874.730 1057.810 ;
        RECT 875.570 1056.750 1041.800 1057.810 ;
        RECT 15.740 4.280 1041.800 1056.750 ;
        RECT 15.740 4.000 74.790 4.280 ;
        RECT 75.630 4.000 224.750 4.280 ;
        RECT 225.590 4.000 374.710 4.280 ;
        RECT 375.550 4.000 524.670 4.280 ;
        RECT 525.510 4.000 674.630 4.280 ;
        RECT 675.470 4.000 824.590 4.280 ;
        RECT 825.430 4.000 974.550 4.280 ;
        RECT 975.390 4.000 1041.800 4.280 ;
      LAYER met3 ;
        RECT 21.040 10.715 1041.600 1050.085 ;
      LAYER met4 ;
        RECT 63.775 11.735 97.440 1039.545 ;
        RECT 99.840 11.735 174.240 1039.545 ;
        RECT 176.640 11.735 251.040 1039.545 ;
        RECT 253.440 11.735 327.840 1039.545 ;
        RECT 330.240 11.735 404.640 1039.545 ;
        RECT 407.040 11.735 481.440 1039.545 ;
        RECT 483.840 11.735 558.240 1039.545 ;
        RECT 560.640 11.735 635.040 1039.545 ;
        RECT 637.440 11.735 711.840 1039.545 ;
        RECT 714.240 11.735 788.640 1039.545 ;
        RECT 791.040 11.735 865.440 1039.545 ;
        RECT 867.840 11.735 942.240 1039.545 ;
        RECT 944.640 11.735 1019.040 1039.545 ;
        RECT 1021.440 11.735 1041.145 1039.545 ;
  END
END user_proj_example
END LIBRARY

