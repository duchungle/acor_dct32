VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN iClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.350 3517.600 2433.910 3524.800 ;
    END
  END iClk
  PIN iRst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 292.820 2924.800 294.020 ;
    END
  END iRst_n
  PIN iSDAT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.990 3517.600 1460.550 3524.800 ;
    END
  END iSDAT
  PIN iSVAL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1759.580 2.400 1760.780 ;
    END
  END iSVAL
  PIN iSize[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2638.820 2924.800 2640.020 ;
    END
  END iSize[0]
  PIN iSize[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.630 3517.600 487.190 3524.800 ;
    END
  END iSize[1]
  PIN iSize[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3225.660 2924.800 3226.860 ;
    END
  END iSize[2]
  PIN iValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 878.980 2924.800 880.180 ;
    END
  END iValid
  PIN oSDAT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1465.820 2924.800 1467.020 ;
    END
  END oSDAT
  PIN oSVAL
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2052.660 2924.800 2053.860 ;
    END
  END oSVAL
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.330 2934.450 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 194.330 2934.450 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 374.330 2934.450 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 554.330 2934.450 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 734.330 2934.450 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 914.330 2934.450 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1094.330 2934.450 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1274.330 2934.450 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1454.330 2934.450 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1634.330 2934.450 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1814.330 2934.450 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1994.330 2934.450 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2174.330 2934.450 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2354.330 2934.450 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2534.330 2934.450 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2714.330 2934.450 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2894.330 2934.450 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3074.330 2934.450 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3254.330 2934.450 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3434.330 2934.450 3437.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -9.470 912.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 -9.470 1092.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -9.470 1272.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 -9.470 1452.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 -9.470 1632.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -9.470 1812.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 -9.470 192.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 -9.470 372.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 -9.470 552.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 -9.470 732.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 2061.030 912.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 2061.030 1092.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 2061.030 1272.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 2061.030 1452.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 2061.030 1632.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 2061.030 1812.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 -9.470 1992.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 -9.470 2172.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 -9.470 2352.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -9.470 2532.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -9.470 2712.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 -9.470 2892.070 3529.150 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 32.930 2944.050 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 212.930 2944.050 216.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 392.930 2944.050 396.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 572.930 2944.050 576.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 752.930 2944.050 756.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 932.930 2944.050 936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1112.930 2944.050 1116.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1292.930 2944.050 1296.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1472.930 2944.050 1476.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1652.930 2944.050 1656.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1832.930 2944.050 1836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2012.930 2944.050 2016.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2192.930 2944.050 2196.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2372.930 2944.050 2376.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2552.930 2944.050 2556.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2732.930 2944.050 2736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2912.930 2944.050 2916.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3092.930 2944.050 3096.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3272.930 2944.050 3276.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3452.930 2944.050 3456.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 -19.070 930.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 -19.070 1110.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 -19.070 1290.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 -19.070 1470.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 -19.070 1650.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 -19.070 1830.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -19.070 30.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 -19.070 210.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 -19.070 390.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 -19.070 570.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 -19.070 750.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 2061.030 930.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 2061.030 1110.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 2061.030 1290.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 2061.030 1470.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 2061.030 1650.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 2061.030 1830.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 -19.070 2010.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 -19.070 2190.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 -19.070 2370.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 -19.070 2550.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 -19.070 2730.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.570 -19.070 2910.670 3538.750 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 51.530 2953.650 54.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 231.530 2953.650 234.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 411.530 2953.650 414.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 591.530 2953.650 594.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 771.530 2953.650 774.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 951.530 2953.650 954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1131.530 2953.650 1134.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1311.530 2953.650 1314.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1491.530 2953.650 1494.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1671.530 2953.650 1674.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1851.530 2953.650 1854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2031.530 2953.650 2034.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2211.530 2953.650 2214.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2391.530 2953.650 2394.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2571.530 2953.650 2574.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2751.530 2953.650 2754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2931.530 2953.650 2934.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3111.530 2953.650 3114.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3291.530 2953.650 3294.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3471.530 2953.650 3474.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 -28.670 949.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 -28.670 1129.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 -28.670 1309.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 -28.670 1489.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 -28.670 1669.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 -28.670 1849.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 -28.670 49.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 -28.670 229.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 -28.670 409.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 -28.670 589.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 -28.670 769.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 2061.030 949.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 2061.030 1129.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 2061.030 1309.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 2061.030 1489.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 2061.030 1669.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 2061.030 1849.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 -28.670 2029.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 -28.670 2209.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 -28.670 2389.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 -28.670 2569.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 -28.670 2749.270 3548.350 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 250.130 2963.250 253.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 430.130 2963.250 433.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 610.130 2963.250 613.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 790.130 2963.250 793.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 970.130 2963.250 973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 -38.270 967.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 -38.270 1147.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 -38.270 1327.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 -38.270 1507.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 -38.270 1687.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 -38.270 1867.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 -38.270 247.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 -38.270 427.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 -38.270 607.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 -38.270 787.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 2061.030 967.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 2061.030 1147.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 2061.030 1327.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 2061.030 1507.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 2061.030 1687.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 2061.030 1867.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 -38.270 2047.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 -38.270 2227.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 -38.270 2407.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 -38.270 2587.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 -38.270 2767.870 3557.950 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 141.530 2953.650 144.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 321.530 2953.650 324.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 501.530 2953.650 504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 681.530 2953.650 684.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 861.530 2953.650 864.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1041.530 2953.650 1044.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1221.530 2953.650 1224.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1401.530 2953.650 1404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1581.530 2953.650 1584.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1761.530 2953.650 1764.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1941.530 2953.650 1944.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2121.530 2953.650 2124.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2301.530 2953.650 2304.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2481.530 2953.650 2484.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2661.530 2953.650 2664.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2841.530 2953.650 2844.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3021.530 2953.650 3024.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3381.530 2953.650 3384.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1036.170 -28.670 1039.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 -28.670 1219.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 -28.670 1399.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 -28.670 1579.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 -28.670 1759.270 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.170 -28.670 139.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 -28.670 319.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 -28.670 499.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 -28.670 679.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 -28.670 859.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1036.170 2061.030 1039.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 2061.030 1219.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 2061.030 1399.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 2061.030 1579.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 2061.030 1759.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 -28.670 1939.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 -28.670 2119.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 -28.670 2299.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 -28.670 2479.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2656.170 -28.670 2659.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.170 -28.670 2839.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 160.130 2963.250 163.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 340.130 2963.250 343.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 520.130 2963.250 523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 700.130 2963.250 703.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 880.130 2963.250 883.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1060.130 2963.250 1063.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1240.130 2963.250 1243.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1420.130 2963.250 1423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1600.130 2963.250 1603.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1780.130 2963.250 1783.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1960.130 2963.250 1963.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2140.130 2963.250 2143.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2320.130 2963.250 2323.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2500.130 2963.250 2503.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2680.130 2963.250 2683.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2860.130 2963.250 2863.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3040.130 2963.250 3043.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3400.130 2963.250 3403.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 -38.270 877.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.770 -38.270 1057.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 -38.270 1237.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 -38.270 1417.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 -38.270 1597.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 -38.270 1777.870 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.770 -38.270 157.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 -38.270 337.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 -38.270 517.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 -38.270 697.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 2061.030 877.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.770 2061.030 1057.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 2061.030 1237.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 2061.030 1417.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 2061.030 1597.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 2061.030 1777.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 -38.270 1957.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 -38.270 2137.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 -38.270 2317.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 -38.270 2497.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2674.770 -38.270 2677.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.770 -38.270 2857.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 104.330 2934.450 107.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 284.330 2934.450 287.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 464.330 2934.450 467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 644.330 2934.450 647.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 824.330 2934.450 827.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1004.330 2934.450 1007.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1184.330 2934.450 1187.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1364.330 2934.450 1367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1544.330 2934.450 1547.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1724.330 2934.450 1727.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1904.330 2934.450 1907.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2084.330 2934.450 2087.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2264.330 2934.450 2267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2444.330 2934.450 2447.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2624.330 2934.450 2627.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2804.330 2934.450 2807.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2984.330 2934.450 2987.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3164.330 2934.450 3167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3344.330 2934.450 3347.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 -9.470 1002.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 -9.470 1182.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 -9.470 1362.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 -9.470 1542.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 -9.470 1722.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 -9.470 1902.070 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 -9.470 102.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 -9.470 282.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 -9.470 462.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 -9.470 642.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 -9.470 822.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 2061.030 1002.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 2061.030 1182.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 2061.030 1362.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 2061.030 1542.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 2061.030 1722.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 2061.030 1902.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 -9.470 2082.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 -9.470 2262.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 -9.470 2442.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 -9.470 2622.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 -9.470 2802.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 122.930 2944.050 126.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 302.930 2944.050 306.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 482.930 2944.050 486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 662.930 2944.050 666.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 842.930 2944.050 846.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1022.930 2944.050 1026.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1202.930 2944.050 1206.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1382.930 2944.050 1386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1562.930 2944.050 1566.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1742.930 2944.050 1746.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1922.930 2944.050 1926.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2102.930 2944.050 2106.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2282.930 2944.050 2286.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2462.930 2944.050 2466.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2642.930 2944.050 2646.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2822.930 2944.050 2826.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3002.930 2944.050 3006.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3362.930 2944.050 3366.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.570 -19.070 1020.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 -19.070 1200.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 -19.070 1380.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 -19.070 1560.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 -19.070 1740.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 -19.070 1920.670 980.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.570 -19.070 120.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 -19.070 300.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 -19.070 480.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 -19.070 660.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 -19.070 840.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.570 2061.030 1020.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 2061.030 1200.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 2061.030 1380.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 2061.030 1560.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 2061.030 1740.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 2061.030 1920.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 -19.070 2100.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 -19.070 2280.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 -19.070 2460.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.570 -19.070 2640.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.570 -19.070 2820.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 880.520 1000.795 1919.660 2040.005 ;
      LAYER met1 ;
        RECT 17.090 296.520 2901.150 3501.620 ;
      LAYER met2 ;
        RECT 17.110 3517.320 486.350 3518.050 ;
        RECT 487.470 3517.320 1459.710 3518.050 ;
        RECT 1460.830 3517.320 2433.070 3518.050 ;
        RECT 2434.190 3517.320 2901.130 3518.050 ;
        RECT 17.110 293.235 2901.130 3517.320 ;
      LAYER met3 ;
        RECT 2.400 3225.260 2917.200 3226.425 ;
        RECT 2.400 2640.420 2917.600 3225.260 ;
        RECT 2.400 2638.420 2917.200 2640.420 ;
        RECT 2.400 2054.260 2917.600 2638.420 ;
        RECT 2.400 2052.260 2917.200 2054.260 ;
        RECT 2.400 1761.180 2917.600 2052.260 ;
        RECT 2.800 1759.180 2917.600 1761.180 ;
        RECT 2.400 1467.420 2917.600 1759.180 ;
        RECT 2.400 1465.420 2917.200 1467.420 ;
        RECT 2.400 880.580 2917.600 1465.420 ;
        RECT 2.400 878.580 2917.200 880.580 ;
        RECT 2.400 294.420 2917.600 878.580 ;
        RECT 2.400 293.255 2917.200 294.420 ;
      LAYER met4 ;
        RECT 896.040 1000.640 1916.145 2040.160 ;
  END
END user_project_wrapper
END LIBRARY

