magic
tech sky130A
magscale 1 2
timestamp 1654564264
<< obsli1 >>
rect 176104 200159 383932 408001
<< obsm1 >>
rect 3418 59304 580230 700324
<< metal2 >>
rect 97326 703520 97438 704960
rect 291998 703520 292110 704960
rect 486670 703520 486782 704960
<< obsm2 >>
rect 3422 703464 97270 703610
rect 97494 703464 291942 703610
rect 292166 703464 486614 703610
rect 486838 703464 580226 703610
rect 3422 58647 580226 703464
<< metal3 >>
rect 583520 645132 584960 645372
rect 583520 527764 584960 528004
rect 583520 410532 584960 410772
rect -960 351916 480 352156
rect 583520 293164 584960 293404
rect 583520 175796 584960 176036
rect 583520 58564 584960 58804
<< obsm3 >>
rect 480 645052 583440 645285
rect 480 528084 583520 645052
rect 480 527684 583440 528084
rect 480 410852 583520 527684
rect 480 410452 583440 410852
rect 480 352236 583520 410452
rect 560 351836 583520 352236
rect 480 293484 583520 351836
rect 480 293084 583440 293484
rect 480 176116 583520 293084
rect 480 175716 583440 176116
rect 480 58884 583520 175716
rect 480 58651 583440 58884
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 9234 -5734 9854 709670
rect 12954 -7654 13574 711590
rect 19794 -1894 20414 705830
rect 23514 -3814 24134 707750
rect 27234 -5734 27854 709670
rect 30954 -7654 31574 711590
rect 37794 -1894 38414 705830
rect 41514 -3814 42134 707750
rect 45234 -5734 45854 709670
rect 48954 -7654 49574 711590
rect 55794 -1894 56414 705830
rect 59514 -3814 60134 707750
rect 63234 -5734 63854 709670
rect 66954 -7654 67574 711590
rect 73794 -1894 74414 705830
rect 77514 -3814 78134 707750
rect 81234 -5734 81854 709670
rect 84954 -7654 85574 711590
rect 91794 -1894 92414 705830
rect 95514 -3814 96134 707750
rect 99234 -5734 99854 709670
rect 102954 -7654 103574 711590
rect 109794 -1894 110414 705830
rect 113514 -3814 114134 707750
rect 117234 -5734 117854 709670
rect 120954 -7654 121574 711590
rect 127794 -1894 128414 705830
rect 131514 -3814 132134 707750
rect 135234 -5734 135854 709670
rect 138954 -7654 139574 711590
rect 145794 -1894 146414 705830
rect 149514 -3814 150134 707750
rect 153234 -5734 153854 709670
rect 156954 -7654 157574 711590
rect 163794 -1894 164414 705830
rect 167514 -3814 168134 707750
rect 171234 -5734 171854 709670
rect 174954 412206 175574 711590
rect 181794 412206 182414 705830
rect 185514 412206 186134 707750
rect 189234 412206 189854 709670
rect 192954 412206 193574 711590
rect 199794 412206 200414 705830
rect 203514 412206 204134 707750
rect 207234 412206 207854 709670
rect 210954 412206 211574 711590
rect 217794 412206 218414 705830
rect 221514 412206 222134 707750
rect 225234 412206 225854 709670
rect 228954 412206 229574 711590
rect 235794 412206 236414 705830
rect 239514 412206 240134 707750
rect 243234 412206 243854 709670
rect 246954 412206 247574 711590
rect 253794 412206 254414 705830
rect 257514 412206 258134 707750
rect 261234 412206 261854 709670
rect 264954 412206 265574 711590
rect 271794 412206 272414 705830
rect 275514 412206 276134 707750
rect 279234 412206 279854 709670
rect 282954 412206 283574 711590
rect 289794 412206 290414 705830
rect 293514 412206 294134 707750
rect 297234 412206 297854 709670
rect 300954 412206 301574 711590
rect 307794 412206 308414 705830
rect 311514 412206 312134 707750
rect 315234 412206 315854 709670
rect 318954 412206 319574 711590
rect 325794 412206 326414 705830
rect 329514 412206 330134 707750
rect 333234 412206 333854 709670
rect 336954 412206 337574 711590
rect 343794 412206 344414 705830
rect 347514 412206 348134 707750
rect 351234 412206 351854 709670
rect 354954 412206 355574 711590
rect 361794 412206 362414 705830
rect 365514 412206 366134 707750
rect 369234 412206 369854 709670
rect 372954 412206 373574 711590
rect 379794 412206 380414 705830
rect 383514 412206 384134 707750
rect 174954 -7654 175574 196000
rect 181794 -1894 182414 196000
rect 185514 -3814 186134 196000
rect 189234 -5734 189854 196000
rect 192954 -7654 193574 196000
rect 199794 -1894 200414 196000
rect 203514 -3814 204134 196000
rect 207234 -5734 207854 196000
rect 210954 -7654 211574 196000
rect 217794 -1894 218414 196000
rect 221514 -3814 222134 196000
rect 225234 -5734 225854 196000
rect 228954 -7654 229574 196000
rect 235794 -1894 236414 196000
rect 239514 -3814 240134 196000
rect 243234 -5734 243854 196000
rect 246954 -7654 247574 196000
rect 253794 -1894 254414 196000
rect 257514 -3814 258134 196000
rect 261234 -5734 261854 196000
rect 264954 -7654 265574 196000
rect 271794 -1894 272414 196000
rect 275514 -3814 276134 196000
rect 279234 -5734 279854 196000
rect 282954 -7654 283574 196000
rect 289794 -1894 290414 196000
rect 293514 -3814 294134 196000
rect 297234 -5734 297854 196000
rect 300954 -7654 301574 196000
rect 307794 -1894 308414 196000
rect 311514 -3814 312134 196000
rect 315234 -5734 315854 196000
rect 318954 -7654 319574 196000
rect 325794 -1894 326414 196000
rect 329514 -3814 330134 196000
rect 333234 -5734 333854 196000
rect 336954 -7654 337574 196000
rect 343794 -1894 344414 196000
rect 347514 -3814 348134 196000
rect 351234 -5734 351854 196000
rect 354954 -7654 355574 196000
rect 361794 -1894 362414 196000
rect 365514 -3814 366134 196000
rect 369234 -5734 369854 196000
rect 372954 -7654 373574 196000
rect 379794 -1894 380414 196000
rect 383514 -3814 384134 196000
rect 387234 -5734 387854 709670
rect 390954 -7654 391574 711590
rect 397794 -1894 398414 705830
rect 401514 -3814 402134 707750
rect 405234 -5734 405854 709670
rect 408954 -7654 409574 711590
rect 415794 -1894 416414 705830
rect 419514 -3814 420134 707750
rect 423234 -5734 423854 709670
rect 426954 -7654 427574 711590
rect 433794 -1894 434414 705830
rect 437514 -3814 438134 707750
rect 441234 -5734 441854 709670
rect 444954 -7654 445574 711590
rect 451794 -1894 452414 705830
rect 455514 -3814 456134 707750
rect 459234 -5734 459854 709670
rect 462954 -7654 463574 711590
rect 469794 -1894 470414 705830
rect 473514 -3814 474134 707750
rect 477234 -5734 477854 709670
rect 480954 -7654 481574 711590
rect 487794 -1894 488414 705830
rect 491514 -3814 492134 707750
rect 495234 -5734 495854 709670
rect 498954 -7654 499574 711590
rect 505794 -1894 506414 705830
rect 509514 -3814 510134 707750
rect 513234 -5734 513854 709670
rect 516954 -7654 517574 711590
rect 523794 -1894 524414 705830
rect 527514 -3814 528134 707750
rect 531234 -5734 531854 709670
rect 534954 -7654 535574 711590
rect 541794 -1894 542414 705830
rect 545514 -3814 546134 707750
rect 549234 -5734 549854 709670
rect 552954 -7654 553574 711590
rect 559794 -1894 560414 705830
rect 563514 -3814 564134 707750
rect 567234 -5734 567854 709670
rect 570954 -7654 571574 711590
rect 577794 -1894 578414 705830
rect 581514 -3814 582134 707750
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 179208 200128 383229 408032
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -6806 694306 590730 694926
rect -4886 690586 588810 691206
rect -2966 686866 586890 687486
rect -8726 680026 592650 680646
rect -6806 676306 590730 676926
rect -4886 672586 588810 673206
rect -2966 668866 586890 669486
rect -8726 662026 592650 662646
rect -6806 658306 590730 658926
rect -4886 654586 588810 655206
rect -2966 650866 586890 651486
rect -8726 644026 592650 644646
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -2966 632866 586890 633486
rect -8726 626026 592650 626646
rect -6806 622306 590730 622926
rect -4886 618586 588810 619206
rect -2966 614866 586890 615486
rect -8726 608026 592650 608646
rect -6806 604306 590730 604926
rect -4886 600586 588810 601206
rect -2966 596866 586890 597486
rect -8726 590026 592650 590646
rect -6806 586306 590730 586926
rect -4886 582586 588810 583206
rect -2966 578866 586890 579486
rect -8726 572026 592650 572646
rect -6806 568306 590730 568926
rect -4886 564586 588810 565206
rect -2966 560866 586890 561486
rect -8726 554026 592650 554646
rect -6806 550306 590730 550926
rect -4886 546586 588810 547206
rect -2966 542866 586890 543486
rect -8726 536026 592650 536646
rect -6806 532306 590730 532926
rect -4886 528586 588810 529206
rect -2966 524866 586890 525486
rect -8726 518026 592650 518646
rect -6806 514306 590730 514926
rect -4886 510586 588810 511206
rect -2966 506866 586890 507486
rect -8726 500026 592650 500646
rect -6806 496306 590730 496926
rect -4886 492586 588810 493206
rect -2966 488866 586890 489486
rect -8726 482026 592650 482646
rect -6806 478306 590730 478926
rect -4886 474586 588810 475206
rect -2966 470866 586890 471486
rect -8726 464026 592650 464646
rect -6806 460306 590730 460926
rect -4886 456586 588810 457206
rect -2966 452866 586890 453486
rect -8726 446026 592650 446646
rect -6806 442306 590730 442926
rect -4886 438586 588810 439206
rect -2966 434866 586890 435486
rect -8726 428026 592650 428646
rect -6806 424306 590730 424926
rect -4886 420586 588810 421206
rect -2966 416866 586890 417486
rect -8726 410026 592650 410646
rect -6806 406306 590730 406926
rect -4886 402586 588810 403206
rect -2966 398866 586890 399486
rect -8726 392026 592650 392646
rect -6806 388306 590730 388926
rect -4886 384586 588810 385206
rect -2966 380866 586890 381486
rect -8726 374026 592650 374646
rect -6806 370306 590730 370926
rect -4886 366586 588810 367206
rect -2966 362866 586890 363486
rect -8726 356026 592650 356646
rect -6806 352306 590730 352926
rect -4886 348586 588810 349206
rect -2966 344866 586890 345486
rect -8726 338026 592650 338646
rect -6806 334306 590730 334926
rect -4886 330586 588810 331206
rect -2966 326866 586890 327486
rect -8726 320026 592650 320646
rect -6806 316306 590730 316926
rect -4886 312586 588810 313206
rect -2966 308866 586890 309486
rect -8726 302026 592650 302646
rect -6806 298306 590730 298926
rect -4886 294586 588810 295206
rect -2966 290866 586890 291486
rect -8726 284026 592650 284646
rect -6806 280306 590730 280926
rect -4886 276586 588810 277206
rect -2966 272866 586890 273486
rect -8726 266026 592650 266646
rect -6806 262306 590730 262926
rect -4886 258586 588810 259206
rect -2966 254866 586890 255486
rect -8726 248026 592650 248646
rect -6806 244306 590730 244926
rect -4886 240586 588810 241206
rect -2966 236866 586890 237486
rect -8726 230026 592650 230646
rect -6806 226306 590730 226926
rect -4886 222586 588810 223206
rect -2966 218866 586890 219486
rect -8726 212026 592650 212646
rect -6806 208306 590730 208926
rect -4886 204586 588810 205206
rect -2966 200866 586890 201486
rect -8726 194026 592650 194646
rect -6806 190306 590730 190926
rect -4886 186586 588810 187206
rect -2966 182866 586890 183486
rect -8726 176026 592650 176646
rect -6806 172306 590730 172926
rect -4886 168586 588810 169206
rect -2966 164866 586890 165486
rect -8726 158026 592650 158646
rect -6806 154306 590730 154926
rect -4886 150586 588810 151206
rect -2966 146866 586890 147486
rect -8726 140026 592650 140646
rect -6806 136306 590730 136926
rect -4886 132586 588810 133206
rect -2966 128866 586890 129486
rect -8726 122026 592650 122646
rect -6806 118306 590730 118926
rect -4886 114586 588810 115206
rect -2966 110866 586890 111486
rect -8726 104026 592650 104646
rect -6806 100306 590730 100926
rect -4886 96586 588810 97206
rect -2966 92866 586890 93486
rect -8726 86026 592650 86646
rect -6806 82306 590730 82926
rect -4886 78586 588810 79206
rect -2966 74866 586890 75486
rect -8726 68026 592650 68646
rect -6806 64306 590730 64926
rect -4886 60586 588810 61206
rect -2966 56866 586890 57486
rect -8726 50026 592650 50646
rect -6806 46306 590730 46926
rect -4886 42586 588810 43206
rect -2966 38866 586890 39486
rect -8726 32026 592650 32646
rect -6806 28306 590730 28926
rect -4886 24586 588810 25206
rect -2966 20866 586890 21486
rect -8726 14026 592650 14646
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal2 s 486670 703520 486782 704960 6 iClk
port 1 nsew signal input
rlabel metal3 s 583520 58564 584960 58804 6 iRst_n
port 2 nsew signal input
rlabel metal2 s 291998 703520 292110 704960 6 iSDAT
port 3 nsew signal input
rlabel metal3 s -960 351916 480 352156 4 iSVAL
port 4 nsew signal input
rlabel metal3 s 583520 527764 584960 528004 6 iSize[0]
port 5 nsew signal input
rlabel metal2 s 97326 703520 97438 704960 6 iSize[1]
port 6 nsew signal input
rlabel metal3 s 583520 645132 584960 645372 6 iSize[2]
port 7 nsew signal input
rlabel metal3 s 583520 175796 584960 176036 6 iValid
port 8 nsew signal input
rlabel metal3 s 583520 293164 584960 293404 6 oSDAT
port 9 nsew signal output
rlabel metal3 s 583520 410532 584960 410772 6 oSVAL
port 10 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 11 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 11 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 11 nsew power input
rlabel metal4 s 181794 -1894 182414 196000 6 vccd1
port 11 nsew power input
rlabel metal4 s 217794 -1894 218414 196000 6 vccd1
port 11 nsew power input
rlabel metal4 s 253794 -1894 254414 196000 6 vccd1
port 11 nsew power input
rlabel metal4 s 289794 -1894 290414 196000 6 vccd1
port 11 nsew power input
rlabel metal4 s 325794 -1894 326414 196000 6 vccd1
port 11 nsew power input
rlabel metal4 s 361794 -1894 362414 196000 6 vccd1
port 11 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 11 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 11 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 181794 412206 182414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 217794 412206 218414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 253794 412206 254414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 289794 412206 290414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 325794 412206 326414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 361794 412206 362414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 11 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 11 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 12 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 12 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 12 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 12 nsew power input
rlabel metal4 s 185514 -3814 186134 196000 6 vccd2
port 12 nsew power input
rlabel metal4 s 221514 -3814 222134 196000 6 vccd2
port 12 nsew power input
rlabel metal4 s 257514 -3814 258134 196000 6 vccd2
port 12 nsew power input
rlabel metal4 s 293514 -3814 294134 196000 6 vccd2
port 12 nsew power input
rlabel metal4 s 329514 -3814 330134 196000 6 vccd2
port 12 nsew power input
rlabel metal4 s 365514 -3814 366134 196000 6 vccd2
port 12 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 12 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 12 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 185514 412206 186134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 221514 412206 222134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 257514 412206 258134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 293514 412206 294134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 329514 412206 330134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 365514 412206 366134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 12 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 12 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 13 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 13 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 13 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 13 nsew power input
rlabel metal4 s 189234 -5734 189854 196000 6 vdda1
port 13 nsew power input
rlabel metal4 s 225234 -5734 225854 196000 6 vdda1
port 13 nsew power input
rlabel metal4 s 261234 -5734 261854 196000 6 vdda1
port 13 nsew power input
rlabel metal4 s 297234 -5734 297854 196000 6 vdda1
port 13 nsew power input
rlabel metal4 s 333234 -5734 333854 196000 6 vdda1
port 13 nsew power input
rlabel metal4 s 369234 -5734 369854 196000 6 vdda1
port 13 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 13 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 13 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 189234 412206 189854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 225234 412206 225854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 261234 412206 261854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 297234 412206 297854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 333234 412206 333854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 369234 412206 369854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 13 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 13 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 14 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 14 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 14 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 14 nsew power input
rlabel metal4 s 192954 -7654 193574 196000 6 vdda2
port 14 nsew power input
rlabel metal4 s 228954 -7654 229574 196000 6 vdda2
port 14 nsew power input
rlabel metal4 s 264954 -7654 265574 196000 6 vdda2
port 14 nsew power input
rlabel metal4 s 300954 -7654 301574 196000 6 vdda2
port 14 nsew power input
rlabel metal4 s 336954 -7654 337574 196000 6 vdda2
port 14 nsew power input
rlabel metal4 s 372954 -7654 373574 196000 6 vdda2
port 14 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 14 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 14 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 192954 412206 193574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 228954 412206 229574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 264954 412206 265574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 300954 412206 301574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 336954 412206 337574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 372954 412206 373574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 14 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 14 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 15 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 207234 -5734 207854 196000 6 vssa1
port 15 nsew ground input
rlabel metal4 s 243234 -5734 243854 196000 6 vssa1
port 15 nsew ground input
rlabel metal4 s 279234 -5734 279854 196000 6 vssa1
port 15 nsew ground input
rlabel metal4 s 315234 -5734 315854 196000 6 vssa1
port 15 nsew ground input
rlabel metal4 s 351234 -5734 351854 196000 6 vssa1
port 15 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 15 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 207234 412206 207854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 243234 412206 243854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 279234 412206 279854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 315234 412206 315854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 351234 412206 351854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 15 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 15 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 16 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 174954 -7654 175574 196000 6 vssa2
port 16 nsew ground input
rlabel metal4 s 210954 -7654 211574 196000 6 vssa2
port 16 nsew ground input
rlabel metal4 s 246954 -7654 247574 196000 6 vssa2
port 16 nsew ground input
rlabel metal4 s 282954 -7654 283574 196000 6 vssa2
port 16 nsew ground input
rlabel metal4 s 318954 -7654 319574 196000 6 vssa2
port 16 nsew ground input
rlabel metal4 s 354954 -7654 355574 196000 6 vssa2
port 16 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 16 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 174954 412206 175574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 210954 412206 211574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 246954 412206 247574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 282954 412206 283574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 318954 412206 319574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 354954 412206 355574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 16 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 16 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 17 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 199794 -1894 200414 196000 6 vssd1
port 17 nsew ground input
rlabel metal4 s 235794 -1894 236414 196000 6 vssd1
port 17 nsew ground input
rlabel metal4 s 271794 -1894 272414 196000 6 vssd1
port 17 nsew ground input
rlabel metal4 s 307794 -1894 308414 196000 6 vssd1
port 17 nsew ground input
rlabel metal4 s 343794 -1894 344414 196000 6 vssd1
port 17 nsew ground input
rlabel metal4 s 379794 -1894 380414 196000 6 vssd1
port 17 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 17 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 199794 412206 200414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 235794 412206 236414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 271794 412206 272414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 307794 412206 308414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 343794 412206 344414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 379794 412206 380414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 17 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 17 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 18 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 203514 -3814 204134 196000 6 vssd2
port 18 nsew ground input
rlabel metal4 s 239514 -3814 240134 196000 6 vssd2
port 18 nsew ground input
rlabel metal4 s 275514 -3814 276134 196000 6 vssd2
port 18 nsew ground input
rlabel metal4 s 311514 -3814 312134 196000 6 vssd2
port 18 nsew ground input
rlabel metal4 s 347514 -3814 348134 196000 6 vssd2
port 18 nsew ground input
rlabel metal4 s 383514 -3814 384134 196000 6 vssd2
port 18 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 18 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 203514 412206 204134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 239514 412206 240134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 275514 412206 276134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 311514 412206 312134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 347514 412206 348134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 383514 412206 384134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 18 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 18 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 95772688
string GDS_FILE /home/hung/caravel_mpw6b/caravel_example/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 94941764
<< end >>

