module prince_wrapper (clk,
    encdec,
    next,
    ready,
    reset_n,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    block,
    key,
    result);
 input clk;
 input encdec;
 input next;
 output ready;
 input reset_n;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input [63:0] block;
 input [127:0] key;
 output [63:0] result;


 prince mprj (.clk(clk),
    .encdec(encdec),
    .next(next),
    .ready(ready),
    .reset_n(reset_n),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .block({block[63],
    block[62],
    block[61],
    block[60],
    block[59],
    block[58],
    block[57],
    block[56],
    block[55],
    block[54],
    block[53],
    block[52],
    block[51],
    block[50],
    block[49],
    block[48],
    block[47],
    block[46],
    block[45],
    block[44],
    block[43],
    block[42],
    block[41],
    block[40],
    block[39],
    block[38],
    block[37],
    block[36],
    block[35],
    block[34],
    block[33],
    block[32],
    block[31],
    block[30],
    block[29],
    block[28],
    block[27],
    block[26],
    block[25],
    block[24],
    block[23],
    block[22],
    block[21],
    block[20],
    block[19],
    block[18],
    block[17],
    block[16],
    block[15],
    block[14],
    block[13],
    block[12],
    block[11],
    block[10],
    block[9],
    block[8],
    block[7],
    block[6],
    block[5],
    block[4],
    block[3],
    block[2],
    block[1],
    block[0]}),
    .key({key[127],
    key[126],
    key[125],
    key[124],
    key[123],
    key[122],
    key[121],
    key[120],
    key[119],
    key[118],
    key[117],
    key[116],
    key[115],
    key[114],
    key[113],
    key[112],
    key[111],
    key[110],
    key[109],
    key[108],
    key[107],
    key[106],
    key[105],
    key[104],
    key[103],
    key[102],
    key[101],
    key[100],
    key[99],
    key[98],
    key[97],
    key[96],
    key[95],
    key[94],
    key[93],
    key[92],
    key[91],
    key[90],
    key[89],
    key[88],
    key[87],
    key[86],
    key[85],
    key[84],
    key[83],
    key[82],
    key[81],
    key[80],
    key[79],
    key[78],
    key[77],
    key[76],
    key[75],
    key[74],
    key[73],
    key[72],
    key[71],
    key[70],
    key[69],
    key[68],
    key[67],
    key[66],
    key[65],
    key[64],
    key[63],
    key[62],
    key[61],
    key[60],
    key[59],
    key[58],
    key[57],
    key[56],
    key[55],
    key[54],
    key[53],
    key[52],
    key[51],
    key[50],
    key[49],
    key[48],
    key[47],
    key[46],
    key[45],
    key[44],
    key[43],
    key[42],
    key[41],
    key[40],
    key[39],
    key[38],
    key[37],
    key[36],
    key[35],
    key[34],
    key[33],
    key[32],
    key[31],
    key[30],
    key[29],
    key[28],
    key[27],
    key[26],
    key[25],
    key[24],
    key[23],
    key[22],
    key[21],
    key[20],
    key[19],
    key[18],
    key[17],
    key[16],
    key[15],
    key[14],
    key[13],
    key[12],
    key[11],
    key[10],
    key[9],
    key[8],
    key[7],
    key[6],
    key[5],
    key[4],
    key[3],
    key[2],
    key[1],
    key[0]}),
    .result({result[63],
    result[62],
    result[61],
    result[60],
    result[59],
    result[58],
    result[57],
    result[56],
    result[55],
    result[54],
    result[53],
    result[52],
    result[51],
    result[50],
    result[49],
    result[48],
    result[47],
    result[46],
    result[45],
    result[44],
    result[43],
    result[42],
    result[41],
    result[40],
    result[39],
    result[38],
    result[37],
    result[36],
    result[35],
    result[34],
    result[33],
    result[32],
    result[31],
    result[30],
    result[29],
    result[28],
    result[27],
    result[26],
    result[25],
    result[24],
    result[23],
    result[22],
    result[21],
    result[20],
    result[19],
    result[18],
    result[17],
    result[16],
    result[15],
    result[14],
    result[13],
    result[12],
    result[11],
    result[10],
    result[9],
    result[8],
    result[7],
    result[6],
    result[5],
    result[4],
    result[3],
    result[2],
    result[1],
    result[0]}));
endmodule
