magic
tech sky130A
magscale 1 2
timestamp 1654560687
<< nwell >>
rect 1066 209157 208970 209723
rect 1066 208069 208970 208635
rect 1066 206981 208970 207547
rect 1066 205893 208970 206459
rect 1066 204805 208970 205371
rect 1066 203717 208970 204283
rect 1066 202629 208970 203195
rect 1066 201541 208970 202107
rect 1066 200453 208970 201019
rect 1066 199365 208970 199931
rect 1066 198277 208970 198843
rect 1066 197189 208970 197755
rect 1066 196101 208970 196667
rect 1066 195013 208970 195579
rect 1066 193925 208970 194491
rect 1066 192837 208970 193403
rect 1066 191749 208970 192315
rect 1066 190661 208970 191227
rect 1066 189573 208970 190139
rect 1066 188485 208970 189051
rect 1066 187397 208970 187963
rect 1066 186309 208970 186875
rect 1066 185221 208970 185787
rect 1066 184133 208970 184699
rect 1066 183045 208970 183611
rect 1066 181957 208970 182523
rect 1066 180869 208970 181435
rect 1066 179781 208970 180347
rect 1066 178693 208970 179259
rect 1066 177605 208970 178171
rect 1066 176517 208970 177083
rect 1066 175429 208970 175995
rect 1066 174341 208970 174907
rect 1066 173253 208970 173819
rect 1066 172165 208970 172731
rect 1066 171077 208970 171643
rect 1066 169989 208970 170555
rect 1066 168901 208970 169467
rect 1066 167813 208970 168379
rect 1066 166725 208970 167291
rect 1066 165637 208970 166203
rect 1066 164549 208970 165115
rect 1066 163461 208970 164027
rect 1066 162373 208970 162939
rect 1066 161285 208970 161851
rect 1066 160197 208970 160763
rect 1066 159109 208970 159675
rect 1066 158021 208970 158587
rect 1066 156933 208970 157499
rect 1066 155845 208970 156411
rect 1066 154757 208970 155323
rect 1066 153669 208970 154235
rect 1066 152581 208970 153147
rect 1066 151493 208970 152059
rect 1066 150405 208970 150971
rect 1066 149317 208970 149883
rect 1066 148229 208970 148795
rect 1066 147141 208970 147707
rect 1066 146053 208970 146619
rect 1066 144965 208970 145531
rect 1066 143877 208970 144443
rect 1066 142789 208970 143355
rect 1066 141701 208970 142267
rect 1066 140613 208970 141179
rect 1066 139525 208970 140091
rect 1066 138437 208970 139003
rect 1066 137349 208970 137915
rect 1066 136261 208970 136827
rect 1066 135173 208970 135739
rect 1066 134085 208970 134651
rect 1066 132997 208970 133563
rect 1066 131909 208970 132475
rect 1066 130821 208970 131387
rect 1066 129733 208970 130299
rect 1066 128645 208970 129211
rect 1066 127557 208970 128123
rect 1066 126469 208970 127035
rect 1066 125381 208970 125947
rect 1066 124293 208970 124859
rect 1066 123205 208970 123771
rect 1066 122117 208970 122683
rect 1066 121029 208970 121595
rect 1066 119941 208970 120507
rect 1066 118853 208970 119419
rect 1066 117765 208970 118331
rect 1066 116677 208970 117243
rect 1066 115589 208970 116155
rect 1066 114501 208970 115067
rect 1066 113413 208970 113979
rect 1066 112325 208970 112891
rect 1066 111237 208970 111803
rect 1066 110149 208970 110715
rect 1066 109061 208970 109627
rect 1066 107973 208970 108539
rect 1066 106885 208970 107451
rect 1066 105797 208970 106363
rect 1066 104709 208970 105275
rect 1066 103621 208970 104187
rect 1066 102533 208970 103099
rect 1066 101445 208970 102011
rect 1066 100357 208970 100923
rect 1066 99269 208970 99835
rect 1066 98181 208970 98747
rect 1066 97093 208970 97659
rect 1066 96005 208970 96571
rect 1066 94917 208970 95483
rect 1066 93829 208970 94395
rect 1066 92741 208970 93307
rect 1066 91653 208970 92219
rect 1066 90565 208970 91131
rect 1066 89477 208970 90043
rect 1066 88389 208970 88955
rect 1066 87301 208970 87867
rect 1066 86213 208970 86779
rect 1066 85125 208970 85691
rect 1066 84037 208970 84603
rect 1066 82949 208970 83515
rect 1066 81861 208970 82427
rect 1066 80773 208970 81339
rect 1066 79685 208970 80251
rect 1066 78597 208970 79163
rect 1066 77509 208970 78075
rect 1066 76421 208970 76987
rect 1066 75333 208970 75899
rect 1066 74245 208970 74811
rect 1066 73157 208970 73723
rect 1066 72069 208970 72635
rect 1066 70981 208970 71547
rect 1066 69893 208970 70459
rect 1066 68805 208970 69371
rect 1066 67717 208970 68283
rect 1066 66629 208970 67195
rect 1066 65541 208970 66107
rect 1066 64453 208970 65019
rect 1066 63365 208970 63931
rect 1066 62277 208970 62843
rect 1066 61189 208970 61755
rect 1066 60101 208970 60667
rect 1066 59013 208970 59579
rect 1066 57925 208970 58491
rect 1066 56837 208970 57403
rect 1066 55749 208970 56315
rect 1066 54661 208970 55227
rect 1066 53573 208970 54139
rect 1066 52485 208970 53051
rect 1066 51397 208970 51963
rect 1066 50309 208970 50875
rect 1066 49221 208970 49787
rect 1066 48133 208970 48699
rect 1066 47045 208970 47611
rect 1066 45957 208970 46523
rect 1066 44869 208970 45435
rect 1066 43781 208970 44347
rect 1066 42693 208970 43259
rect 1066 41605 208970 42171
rect 1066 40517 208970 41083
rect 1066 39429 208970 39995
rect 1066 38341 208970 38907
rect 1066 37253 208970 37819
rect 1066 36165 208970 36731
rect 1066 35077 208970 35643
rect 1066 33989 208970 34555
rect 1066 32901 208970 33467
rect 1066 31813 208970 32379
rect 1066 30725 208970 31291
rect 1066 29637 208970 30203
rect 1066 28549 208970 29115
rect 1066 27461 208970 28027
rect 1066 26373 208970 26939
rect 1066 25285 208970 25851
rect 1066 24197 208970 24763
rect 1066 23109 208970 23675
rect 1066 22021 208970 22587
rect 1066 20933 208970 21499
rect 1066 19845 208970 20411
rect 1066 18757 208970 19323
rect 1066 17669 208970 18235
rect 1066 16581 208970 17147
rect 1066 15493 208970 16059
rect 1066 14405 208970 14971
rect 1066 13317 208970 13883
rect 1066 12229 208970 12795
rect 1066 11141 208970 11707
rect 1066 10053 208970 10619
rect 1066 8965 208970 9531
rect 1066 7877 208970 8443
rect 1066 6789 208970 7355
rect 1066 5701 208970 6267
rect 1066 4613 208970 5179
rect 1066 3525 208970 4091
rect 1066 2437 208970 3003
<< obsli1 >>
rect 1104 2159 208932 210001
<< obsm1 >>
rect 1104 2128 208932 210032
<< metal2 >>
rect 34978 211406 35034 212206
rect 104990 211406 105046 212206
rect 175002 211406 175058 212206
rect 15014 0 15070 800
rect 45006 0 45062 800
rect 74998 0 75054 800
rect 104990 0 105046 800
rect 134982 0 135038 800
rect 164974 0 165030 800
rect 194966 0 195022 800
<< obsm2 >>
rect 3148 211350 34922 211562
rect 35090 211350 104934 211562
rect 105102 211350 174946 211562
rect 175114 211350 208360 211562
rect 3148 856 208360 211350
rect 3148 800 14958 856
rect 15126 800 44950 856
rect 45118 800 74942 856
rect 75110 800 104934 856
rect 105102 800 134926 856
rect 135094 800 164918 856
rect 165086 800 194910 856
rect 195078 800 208360 856
<< obsm3 >>
rect 4208 2143 208320 210017
<< metal4 >>
rect 4208 2128 4528 210032
rect 19568 2128 19888 210032
rect 34928 2128 35248 210032
rect 50288 2128 50608 210032
rect 65648 2128 65968 210032
rect 81008 2128 81328 210032
rect 96368 2128 96688 210032
rect 111728 2128 112048 210032
rect 127088 2128 127408 210032
rect 142448 2128 142768 210032
rect 157808 2128 158128 210032
rect 173168 2128 173488 210032
rect 188528 2128 188848 210032
rect 203888 2128 204208 210032
<< obsm4 >>
rect 12755 2347 19488 207909
rect 19968 2347 34848 207909
rect 35328 2347 50208 207909
rect 50688 2347 65568 207909
rect 66048 2347 80928 207909
rect 81408 2347 96288 207909
rect 96768 2347 111648 207909
rect 112128 2347 127008 207909
rect 127488 2347 142368 207909
rect 142848 2347 157728 207909
rect 158208 2347 173088 207909
rect 173568 2347 188448 207909
rect 188928 2347 203808 207909
rect 204288 2347 208229 207909
<< labels >>
rlabel metal2 s 15014 0 15070 800 6 iClk
port 1 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 iRst_n
port 2 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 iSDAT
port 3 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 iSVAL
port 4 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 iSize[0]
port 5 nsew signal input
rlabel metal2 s 175002 211406 175058 212206 6 iSize[1]
port 6 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 iSize[2]
port 7 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 iValid
port 8 nsew signal input
rlabel metal2 s 104990 211406 105046 212206 6 oSDAT
port 9 nsew signal output
rlabel metal2 s 34978 211406 35034 212206 6 oSVAL
port 10 nsew signal output
rlabel metal4 s 4208 2128 4528 210032 6 vccd1
port 11 nsew power input
rlabel metal4 s 34928 2128 35248 210032 6 vccd1
port 11 nsew power input
rlabel metal4 s 65648 2128 65968 210032 6 vccd1
port 11 nsew power input
rlabel metal4 s 96368 2128 96688 210032 6 vccd1
port 11 nsew power input
rlabel metal4 s 127088 2128 127408 210032 6 vccd1
port 11 nsew power input
rlabel metal4 s 157808 2128 158128 210032 6 vccd1
port 11 nsew power input
rlabel metal4 s 188528 2128 188848 210032 6 vccd1
port 11 nsew power input
rlabel metal4 s 19568 2128 19888 210032 6 vssd1
port 12 nsew ground input
rlabel metal4 s 50288 2128 50608 210032 6 vssd1
port 12 nsew ground input
rlabel metal4 s 81008 2128 81328 210032 6 vssd1
port 12 nsew ground input
rlabel metal4 s 111728 2128 112048 210032 6 vssd1
port 12 nsew ground input
rlabel metal4 s 142448 2128 142768 210032 6 vssd1
port 12 nsew ground input
rlabel metal4 s 173168 2128 173488 210032 6 vssd1
port 12 nsew ground input
rlabel metal4 s 203888 2128 204208 210032 6 vssd1
port 12 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 210062 212206
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 94941710
string GDS_FILE /home/hung/caravel_mpw6b/caravel_example/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 1234170
<< end >>

